module top_robotic_arm();

endmodule